// SAP-1 Controller
/*
Controller is the sole independent element of the SAP-1

Controller drives clock and clear signals

Controller drives the enable pins of all other elements
Control logic is driven depending on how designer decodes instructions
into control signals

Controller reads instruction from instruction register as necessary

*/

module SAP_1(instruction, clock, clock_inv, clear, clear_inv, control_word);
  
  input [3:0] instruction;
  input clock;				
  // Clock should be output as a standalone signal generated by controller
  // But since this is verilog implementation, a module cannot generate clock sig and 
  // has to be externally input
  output clock_inv, clear, clear_inv;
  output reg[11:0] control_word;
  
  // these parameters are used to reference control word bits
  parameter Cp = 11;// active high	// program counter count signal
  parameter Ep = 10;// active high	// program counter enable output (to BUS)
  parameter Lm = 9; // active low	// memory address register enable load
  parameter Ce = 8; // active low	// RAM enable output (to BUS)
  parameter Li = 7; // active low	// instruction register load data (from BUS)
  parameter Ei = 6; // active low	// instruction register enable output (to BUS)
  parameter La = 5; // active low	// accumulator load data (from BUS)
  parameter Ea = 4; // active high	// accumulator enable output (to BUS)
  parameter Su = 3; // sub on high	// ALU operation mode
  parameter Eu = 2; // active high	// ALU enable output (to BUS)
  parameter Lb = 1; // active low	// Register B data load (from BUS)
  parameter Lo = 0; // active low	// Output Register data load (from BUS)
  
  reg [5:0] ring_counter;
  reg clear;
  reg [3:0] OP_CODE;
    
  assign clock_inv = ~clock;
  assign clear_inv = ~clear;
  
  // 6 bit ring counter
  always @(negedge clock) begin
    
	if (ring_counter == 6'b000000) begin// system just came alive 
		ring_counter = 6'b000001;
		clear = 1;
	end
	else if (ring_counter == 6'b100000) // completed a full cycle
		ring_counter = 6'b000001;
	else begin
		clear = 0;
		ring_counter = ring_counter * 2;
	end
  end
  
  // Instruction sequence and decoder
  always @(negedge clock) begin

    case (ring_counter)
	  // CON == [Cp Ep Lm' Ce'   Li' Ei' La' Ea   Su Eu Lb' Lo']
    
      // T1 Address State // 1st step of fetch cycle
      6'b000001  : control_word <= 12'b010111100011;
      // Program counter address is transferred to (Ep)
      // Memory address register (Lm')
      
      6'b000010  : control_word <= 12'b101111100011;
      // T2 Increment State // 2nd step of fetch cycle
      // Program counter is set to increment (Cp)
      
      // T3 Memory State // 3rd step of fetch cycle
      6'b000100  : control_word <= 12'b001001100011;
      // RAM instruction is transferred to (Ce')
      // Instruction register (Li')
      
      // T4 State // 1st step of execution cycle
      6'b001000  : begin
		if (instruction == 4'b0000) // LDA routine
			control_word <= 12'b000110100011; // Lm' and Ei' active (low)
		else if (instruction == 4'b0001) //	ADD routine
			control_word <= 12'b000110100011; // Lm' and Ei' active (low)
		else if (instruction == 4'b0010) //	SUB routine
			control_word <= 12'b000110100011; // Lm' and Ei' active (low)
		else if (instruction == 4'b1110) // OUT routine
			control_word <= 12'b001111110010; // Ea and Lo' active
		else if (instruction == 4'b1111) // HLT routine (NOT YET IMPLEMENTED)
			control_word <= 12'b001111100011; // NOP
		else
			control_word <= 12'b001111100011; // NOP
      end
      
      // T5 State // 2nd step of execution cycle
      6'b010000  : begin
		if (instruction == 4'b0000) // LDA routine
			control_word <= 12'b001011000011; // Ce' and La' active (low)
		else if (instruction == 4'b0001) //	ADD routine
			control_word <= 12'b001011100001; // Ce' and Lb' active (low)
		else if (instruction == 4'b0010) //	SUB routine
			control_word <= 12'b001011100001; // Ce' and Lb' active (low)
		else if (instruction == 4'b1110) // OUT routine
			control_word <= 12'b001111100011; // NOP
		else if (instruction == 4'b1111) // HLT routine (NOT YET IMPLEMENTED)
			control_word <= 12'b001111100011; // NOP
		else
			control_word <= 12'b001111100011; // NOP
      end
      
      // T6 State // 3rd step of execution cycle
      6'b100000  : begin
		if (instruction == 4'b0000) // LDA routine
			control_word <= 12'b001111100011; // NOP
		else if (instruction == 4'b0001) //	ADD routine
			control_word <= 12'b000110000111; // Eu and La' active
		else if (instruction == 4'b0010) //	SUB routine
			control_word <= 12'b000110001111; // Eu, Su and La' active
		else if (instruction == 4'b1110) // OUT routine
			control_word <= 12'b001111100011; // NOP
		else if (instruction == 4'b1111) // HLT routine (NOT YET IMPLEMENTED)
			control_word <= 12'b001111100011; // NOP
		else
			control_word <= 12'b001111100011; // NOP	
      end 
      
      default : control_word <= 12'b001111100011; // NOP
    
    endcase
  end
    
endmodule
